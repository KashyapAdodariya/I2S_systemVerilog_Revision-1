`define size 16
`include "i2s_message_logger.sv"
`include "i2s_config.sv"
`include "i2s_coverage.sv"
`include "i2s_transaction.sv"
`include "i2s_interface.sv"
`include "i2s_master_gen.sv"
`include "i2s_master_driver.sv"
`include "i2s_monitor.sv"
`include "i2s_master_agent.sv"
`include "i2s_slave_driver.sv"
`include "i2s_slave_agent.sv"
`include "i2s_scoreboard.sv"
`include "i2s_env.sv"

`ifdef test1
`include "/tests/alteranate_data_stream_mono_left_mode.sv"
`elsif test2
`include "/tests/alteranate_data_stream_mono_right_mode.sv"
`elsif  test3
`include "/tests/alteranate_data_stream_stereo_mode.sv"
`elsif  test4
`include "/tests/change_word_len.sv"
`elsif  test5
`include "/tests/slave_tx_twos_stereo.sv"
`elsif test6
`include "/tests/const_data_stream_mono_left_mode.sv"
`elsif test7
`include "/tests/const_data_stream_mono_right_mode.sv"
`elsif test8
`include "/tests/const_data_stream_stereo_mode.sv"
`elsif test9
`include "/tests/extra_bit_master_tx.sv"
`elsif  test10
`include "/tests/stereo_mode.sv"
`elsif test11
`include "/tests/illegal_word_len.sv"
`elsif  test12
`include "/tests/master_tx_and_slave_rx_wlen_same.sv"
`elsif test13
`include "/tests/master_tx_normal_mono_left.sv"
`elsif test14
`include "/tests/master_tx_normal_mono_right.sv"
`elsif test15
`include "/tests/master_tx_normal_stereo.sv"
`elsif  test16
`include "/tests/master_tx_twos_mono_left.sv"
`elsif test17
`include "/tests/master_tx_twos_mono_right.sv"
`elsif  test18
`include "/tests/master_tx_twos_stereo.sv"
`elsif  test19
`include "/tests/master_tx_wlen_greaterthen_slave_mono_left.sv"
`elsif  test20
`include "/tests/master_tx_wlen_greaterthen_slave_mono_right.sv"
`elsif  test21
`include "/tests/master_tx_wlen_greaterthen_slave_stereo.sv"
`elsif  test22
`include "/tests/mono_left_mode.sv"
`elsif  test23
`include "/tests/mono_right_mode.sv"
`elsif  test24
`include "/tests/rx_word_len_gr_tx_word_len.sv"
`elsif test25
`include "/tests/slave_tx_normal_mono_left.sv"
`elsif  test26
`include "/tests/slave_tx_normal_mono_right.sv"
`elsif  test27
`include "/tests/slave_tx_normal_stereo.sv"
`elsif  test28
`include "/tests/slave_tx_twos_mono_left.sv"
`elsif test29
`include "/tests/slave_tx_twos_mono_right.sv"
`endif


